// Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
// Please do not spread this code without permission 
module mac_array (clk, reset, out_s, in_w, in_n, inst_w, mode, valid);
  parameter act_bw = 2;
  parameter w_bw = 4;
  parameter psum_bw = 16;
  parameter col = 8;
  parameter row = 8;

  input  clk, reset;
  output [2*psum_bw*col-1:0] out_s;
  input  [row*w_bw-1:0] in_w; // inst[1]:execute, inst[0]: kernel loading
  input  [1:0] inst_w;
  input  [2*psum_bw*col-1:0] in_n;
  input mode; //0: 4-bit act and 4-bit weight;    1: 2-bit act and 4-bit weight
  output [col-1:0] valid;


  reg    [2*row-1:0] inst_w_temp;
  wire   [2*psum_bw*col*(row+1)-1:0] temp;
  wire   [row*col-1:0] valid_temp;


  genvar i;
 
  assign out_s = temp[2*psum_bw*col*9-1:2*psum_bw*col*8];
  assign temp[psum_bw*col*1-1:psum_bw*col*0] = 0;
  assign valid = valid_temp[row*col-1:row*col-8];

  for (i=1; i < row+1 ; i=i+1) begin : row_num
      mac_row #(.act_bw(act_bw), .w_bw(w_bw), .psum_bw(psum_bw)) mac_row_instance (
        .clk(clk),
        .reset(reset),
        .mode(mode),
	      .in_w(in_w[w_bw*i-1:w_bw*(i-1)]),
	      .inst_w(inst_w_temp[2*i-1:2*(i-1)]),
	      .in_n(temp[2*psum_bw*col*i-1:2*psum_bw*col*(i-1)]),
        .valid(valid_temp[col*i-1:col*(i-1)]),
	      .out_s(temp[2*psum_bw*col*(i+1)-1:2*psum_bw*col*(i)]));
  end

  always @ (posedge clk) begin

    //valid <= valid_temp[row*col-1:row*col-8];
    // Add new instruction in the lower 2 bits and pass
		// instructions from previous row to the next one
		inst_w_temp <= {inst_w_temp[2*row-3:0], inst_w};

  end

endmodule
